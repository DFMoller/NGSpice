* Electronics 315 - W01L3
* BJT CE with RE gain
* Author: CJ Fourie
* Last mod: 9 February 2021
**************************************

Vs      In     0        0     AC    1     0

VCC     VCC    0        10

RS      in     1        0.5k
R1      VCC    qb       56k
R2      qb     0        12.2k
RC      VCC    out      2k
RE      qe     0        0.4k

CC      1      qb       100m

*       Collector   Base     Emitter   Model
Q1      out         qb       qe        BJT1

.model BJT1 NPN (BF=100 IS=1e-15)

* A zero current source at the output is open during normal simulation
* but is used to measure output resistance later
Io      0      out      ac     0    0

.control
  AC    DEC    1   10k   10k          $  Do ac analysis at single frequency
*  To calculate output resistance, zero the input voltage and apply
*    an ac current at output (if we apply a voltage at the output, it will
*    short the collector to ground - not intended).
  alter @Vs[acmag]=0               $ Set Vs = 0:
  alter @Io[acmag]=1               $ Set Io = 1 A (0 deg phase):
  AC    DEC     1  10k   10k       $ Run AC analysis again
  
  meas ac vi_magn max ac1.v(in) AT=10k    $  Measure ac magnitudes at 10 kHz from first ac analysis
  meas ac ii_magn max ac1.i(vs) AT=10k 
  meas ac vo_magn max ac1.v(out) AT=10k
  meas ac v1_magn max ac1.v(1) AT=10k
  meas ac vo_magn2 max ac2.v(out) AT=10k  $  Measure ac magnitude at 10 kHz from second ac analysis

  let Av = vo_magn/(vi_magn)
  let Ri = v1_magn/(-ii_magn)  
  let Ro = vo_magn2                      $ We know Io[acmag] = 1, so Ro = max(vo_magn2)
  echo
  echo Voltage gain Av = "$&Av" V/V
  echo Input resistance Ri = "$&Ri" Ohm
  echo Closed-loop output resistance Ro = "$&Ro" Ohm
  echo 
.endc
.end