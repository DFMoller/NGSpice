* SPICE model for power amplifier
*-------------------------------------------------------------
* Author: Your Name
* SU student number : 12345679
* Last mod: 21 April 2021
*=============================================================
* Description: This Class-A is used to show (non-)compliance
* specifications and tests for Electronics 315 practical 3
*=============================================================

* YOUR CIRCUIT MUST INCLUDE:
* 1. A voltage source (DC 0) in series with the emitter of Qn, named Vicn, to measure I_{CQn}.
*    Its POSITIVE node must be connected to the emitter of Qn, and named "qne"
*      Example:  Vicn qne nodewhatever  DC  0
* 2. A voltage source (DC 0) in series with the emitter of Qp, named Vicp, to measure I_{CQp}.
*    Its NEGATIVE node must be connected to the emitter of Qp, and named "qpe"
*      Example:  Vicp nodewhateverelse  qpe  DC  0

* Include the transistor models as an external file ("models.cir"); these are standard for the module
.include models.cir

* Define amplifier as a subcircuit to avoid node name clashes in test bench
* subckt name must be "audioamp"
* ---------------------------------------------------------------------------------------------
* Pin sequence must be:  SignalInput+, SpeakerOut+, SpeakerOut-, SupplyVoltage+, SupplyVoltage-
* ---------------------------------------------------------------------------------------------

.subckt  audioamp  in  out  outn  vcc  vee 

* Finally, your circuit is defined below:

* ============== CUT OUT BELOW AND BUILD YOUR CIRCUIT ====================
* Class-B stage - no cross-over support
Q2   VCC    qnb       qne   TIP41C
Vicn qne    noden     DC    0
Q4   VEE    qpb       qpe   TIP41C
Vicp nodep  qpe       DC    0
Q1   VCC    preampout qnb   t2N2219A
Q3   VEE    preampout qpb   t2N2905A
Ren  noden  pwrout    1u
Rep  nodep  pwrout    1u 

*Rbias1  VCC preampof  100
*Rbias2  VEE preampout  100
*Roffset preampof preampout 14

Qpa1   preampout preampin  qpae  t2N2219A
Rbias1 VCC preampin    60k
Rbias2 VEE preampin    80k
Rpac   VCC preampout   200
Rpae   qpae  VEE       50  


Cin  in     preampin  100u
Cout pwrout out       4700u

* ============== CUT OUT ABOVE AND BUILD YOUR CIRCUIT ====================

* low resistance speaker connection to ground (to avoid putting "0" in the .subckt line

Rcable outn 0  1m

.ends
* ============================================


